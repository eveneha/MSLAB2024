ms24.41@localhost.localdomain.14821:1710255337