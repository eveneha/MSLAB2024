package CONSTANTS is
   constant tp_mux : time := 0 ns;
   constant numBit : integer := 64; 
   constant IVDELAY : time := 0.1 ns;
   constant NDDELAY : time := 0.2 ns;
   constant NRDELAY : time := 0.2 ns;
end CONSTANTS;
